`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 20.03.2024 18:05:44
// Design Name: 
// Module Name: mux8to1_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux8to1_tb();
    logic i[7:0],s[2:0],y;
    mux8to1 dut(i[0],i[1],i[2],i[3],i[4],i[5],i[6],i[7],s[0],s[1],s[2],y);
    initial begin
    i = {0,0,0,0,0,0,0,0}; s = {0,0,0}; #20;
    i = {0,0,0,0,0,0,0,1}; s = {0,0,0}; #20;
    i = {0,0,0,0,0,0,0,0}; s = {0,0,1}; #20;
    i = {0,0,0,0,0,0,1,0}; s = {0,0,1}; #20;
    i = {0,0,0,0,0,0,0,0}; s = {0,1,0}; #20;
    i = {0,0,0,0,0,1,0,0}; s = {0,1,0}; #20;
    i = {0,0,0,0,0,0,0,0}; s = {0,1,1}; #20;
    i = {0,0,0,0,1,0,0,0}; s = {0,1,1}; #20;
    i = {0,0,0,0,0,0,0,0}; s = {1,0,0}; #20;
    i = {0,0,0,1,0,0,0,0}; s = {1,0,0}; #20;
    i = {0,0,0,0,0,0,0,0}; s = {1,0,1}; #20;
    i = {0,0,1,0,0,0,0,0}; s = {1,0,1}; #20;
    i = {0,0,0,0,0,0,0,0}; s = {1,1,0}; #20;
    i = {0,1,0,0,0,0,0,0}; s = {1,1,0}; #20;
    i = {0,0,0,0,0,0,0,0}; s = {1,1,1}; #20;
    i = {1,0,0,0,0,0,0,0}; s = {1,1,1}; #20;
    end
endmodule
